.subckt Core_test_flow INM INP OUTM OUTP VBIAS_P VDD VREF VSS
XP1c_0 net020 VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1c_1 net020 VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1c_2 net020 VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1c_3 net020 VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1c_4 net020 VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1c_5 net020 VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1c_6 net020 VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1c_7 net020 VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X20_0 net028 VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X20_1 net028 VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X20_2 net028 VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X20_3 net028 VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X20_4 net028 VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X20_5 net028 VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X20_6 net028 VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X20_7 net028 VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X7_0 vbias_n VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X7_1 vbias_n VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X7_2 vbias_n VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X7_3 vbias_n VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X7_4 vbias_n VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X7_5 vbias_n VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X7_6 vbias_n VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X7_7 vbias_n VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X5_0 VBIAS_P VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X5_1 VBIAS_P VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X5_2 VBIAS_P VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X5_3 VBIAS_P VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X5_4 VBIAS_P VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X5_5 VBIAS_P VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X5_6 VBIAS_P VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X5_7 VBIAS_P VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1a_0 intm VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1a_1 intm VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1a_2 intm VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1a_3 intm VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1a_4 intm VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1a_5 intm VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1a_6 intm VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1a_7 intm VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1a_8 intm VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1a_9 intm VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1a_10 intm VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1a_11 intm VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1a_12 intm VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1a_13 intm VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1a_14 intm VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1a_15 intm VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1a_16 intm VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1a_17 intm VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1a_18 intm VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1a_19 intm VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1b_0 intp VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1b_1 intp VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1b_2 intp VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1b_3 intp VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1b_4 intp VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1b_5 intp VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1b_6 intp VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1b_7 intp VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1b_8 intp VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1b_9 intp VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1b_10 intp VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1b_11 intp VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1b_12 intp VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1b_13 intp VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1b_14 intp VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1b_15 intp VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1b_16 intp VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1b_17 intp VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1b_18 intp VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XP1b_19 intp VBIAS_P VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
XC1_0 net037 OUTM sky130_fd_pr__cap_mim_m3_1 l=5.0e+06u w=5.0e+06u
XC0_0 net047 OUTP sky130_fd_pr__cap_mim_m3_1 l=5.0e+06u w=5.0e+06u
X10_0 net7 vbias_n VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X10_1 net7 vbias_n VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X10_2 net7 vbias_n VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X10_3 net7 vbias_n VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X10_4 net7 vbias_n VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X10_5 net7 vbias_n VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X10_6 net7 vbias_n VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X10_7 net7 vbias_n VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X10_8 net7 vbias_n VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X10_9 net7 vbias_n VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X10_10 net7 vbias_n VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X10_11 net7 vbias_n VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X10_12 net7 vbias_n VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X10_13 net7 vbias_n VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X10_14 net7 vbias_n VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X10_15 net7 vbias_n VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X9_0 OUTM vbias_n VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X9_1 OUTM vbias_n VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X9_2 OUTM vbias_n VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X9_3 OUTM vbias_n VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X9_4 OUTM vbias_n VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X9_5 OUTM vbias_n VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X6_0 OUTP vbias_n VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X6_1 OUTP vbias_n VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X6_2 OUTP vbias_n VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X6_3 OUTP vbias_n VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X6_4 OUTP vbias_n VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X6_5 OUTP vbias_n VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X13_0 vcmfb vcmfb VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X13_1 vcmfb vcmfb VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X12_0 net025 net025 VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X12_1 net025 net025 VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X11_0 net7 vcmfb VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X11_1 net7 vcmfb VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X11_2 net7 vcmfb VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X11_3 net7 vcmfb VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X4_0 vbias_n vbias_n VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X4_1 vbias_n vbias_n VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X4_2 vbias_n vbias_n VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X4_3 vbias_n vbias_n VSS VSS sky130_fd_pr__nfet_01v8_lvt l=2.4e+5u w=2.0e+06u
X19_0 net025 VREF net028 VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X19_1 net025 VREF net028 VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X19_2 net025 VREF net028 VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X19_3 net025 VREF net028 VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X19_4 net025 VREF net028 VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X19_5 net025 VREF net028 VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X19_6 net025 VREF net028 VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X19_7 net025 VREF net028 VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X17_0 net025 VREF net020 VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X17_1 net025 VREF net020 VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X17_2 net025 VREF net020 VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X17_3 net025 VREF net020 VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X17_4 net025 VREF net020 VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X17_5 net025 VREF net020 VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X17_6 net025 VREF net020 VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X17_7 net025 VREF net020 VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X15_0 vcmfb OUTP net020 VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X15_1 vcmfb OUTP net020 VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X15_2 vcmfb OUTP net020 VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X15_3 vcmfb OUTP net020 VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X15_4 vcmfb OUTP net020 VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X15_5 vcmfb OUTP net020 VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X15_6 vcmfb OUTP net020 VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X15_7 vcmfb OUTP net020 VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X25_0 net037 VSS intp VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X25_1 net037 VSS intp VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X25_2 net037 VSS intp VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X25_3 net037 VSS intp VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X25_4 net037 VSS intp VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X25_5 net037 VSS intp VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X25_6 net037 VSS intp VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X25_7 net037 VSS intp VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X25_8 net037 VSS intp VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X25_9 net037 VSS intp VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X25_10 net037 VSS intp VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X25_11 net037 VSS intp VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X23_0 net047 VSS intm VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X23_1 net047 VSS intm VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X23_2 net047 VSS intm VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X23_3 net047 VSS intm VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X23_4 net047 VSS intm VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X23_5 net047 VSS intm VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X23_6 net047 VSS intm VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X23_7 net047 VSS intm VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X23_8 net047 VSS intm VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X23_9 net047 VSS intm VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X23_10 net047 VSS intm VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X23_11 net047 VSS intm VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X3_0 OUTP intm VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X3_1 OUTP intm VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X3_2 OUTP intm VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X3_3 OUTP intm VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X3_4 OUTP intm VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X3_5 OUTP intm VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X3_6 OUTP intm VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X3_7 OUTP intm VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X3_8 OUTP intm VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X3_9 OUTP intm VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X3_10 OUTP intm VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X3_11 OUTP intm VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X1_0 OUTM intp VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X1_1 OUTM intp VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X1_2 OUTM intp VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X1_3 OUTM intp VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X1_4 OUTM intp VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X1_5 OUTM intp VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X1_6 OUTM intp VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X1_7 OUTM intp VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X1_8 OUTM intp VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X1_9 OUTM intp VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X1_10 OUTM intp VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X1_11 OUTM intp VDD VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X18_0 vcmfb OUTM net028 VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X18_1 vcmfb OUTM net028 VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X18_2 vcmfb OUTM net028 VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X18_3 vcmfb OUTM net028 VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X18_4 vcmfb OUTM net028 VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X18_5 vcmfb OUTM net028 VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X18_6 vcmfb OUTM net028 VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X18_7 vcmfb OUTM net028 VDD sky130_fd_pr__pfet_01v8 l=2.4e+5u w=2.0e+06u
X0_0 intp INM net7 VSS sky130_fd_pr__nfet_01v8 l=5.0e+5u w=5.0e+06u
X0_1 intp INM net7 VSS sky130_fd_pr__nfet_01v8 l=5.0e+5u w=5.0e+06u
X0_2 intp INM net7 VSS sky130_fd_pr__nfet_01v8 l=5.0e+5u w=5.0e+06u
X0_3 intp INM net7 VSS sky130_fd_pr__nfet_01v8 l=5.0e+5u w=5.0e+06u
X0_4 intp INM net7 VSS sky130_fd_pr__nfet_01v8 l=5.0e+5u w=5.0e+06u
X0_5 intp INM net7 VSS sky130_fd_pr__nfet_01v8 l=5.0e+5u w=5.0e+06u
X0_6 intp INM net7 VSS sky130_fd_pr__nfet_01v8 l=5.0e+5u w=5.0e+06u
X0_7 intp INM net7 VSS sky130_fd_pr__nfet_01v8 l=5.0e+5u w=5.0e+06u
X0_8 intp INM net7 VSS sky130_fd_pr__nfet_01v8 l=5.0e+5u w=5.0e+06u
X0_9 intp INM net7 VSS sky130_fd_pr__nfet_01v8 l=5.0e+5u w=5.0e+06u
X0_10 intp INM net7 VSS sky130_fd_pr__nfet_01v8 l=5.0e+5u w=5.0e+06u
X0_11 intp INM net7 VSS sky130_fd_pr__nfet_01v8 l=5.0e+5u w=5.0e+06u
X2_0 intm INP net7 VSS sky130_fd_pr__nfet_01v8 l=5.0e+5u w=5.0e+06u
X2_1 intm INP net7 VSS sky130_fd_pr__nfet_01v8 l=5.0e+5u w=5.0e+06u
X2_2 intm INP net7 VSS sky130_fd_pr__nfet_01v8 l=5.0e+5u w=5.0e+06u
X2_3 intm INP net7 VSS sky130_fd_pr__nfet_01v8 l=5.0e+5u w=5.0e+06u
X2_4 intm INP net7 VSS sky130_fd_pr__nfet_01v8 l=5.0e+5u w=5.0e+06u
X2_5 intm INP net7 VSS sky130_fd_pr__nfet_01v8 l=5.0e+5u w=5.0e+06u
X2_6 intm INP net7 VSS sky130_fd_pr__nfet_01v8 l=5.0e+5u w=5.0e+06u
X2_7 intm INP net7 VSS sky130_fd_pr__nfet_01v8 l=5.0e+5u w=5.0e+06u
X2_8 intm INP net7 VSS sky130_fd_pr__nfet_01v8 l=5.0e+5u w=5.0e+06u
X2_9 intm INP net7 VSS sky130_fd_pr__nfet_01v8 l=5.0e+5u w=5.0e+06u
X2_10 intm INP net7 VSS sky130_fd_pr__nfet_01v8 l=5.0e+5u w=5.0e+06u
X2_11 intm INP net7 VSS sky130_fd_pr__nfet_01v8 l=5.0e+5u w=5.0e+06u

.ends
