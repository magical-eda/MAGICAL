.subckt COMPARATOR CLK CROSSN CROSSP GND INTERN INTERP OUTM OUTP VDD VI+ VI-

X0_0 GND INTERN GND GND sky130_fd_pr__nfet_01v8_lvt l=1e+06u w=5.25e+06u 
X22_0 GND INTERP GND GND sky130_fd_pr__nfet_01v8_lvt l=1e+06u w=5.25e+06u
X16_0 OUTM CROSSP GND GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=2.4e+06u
X16_1 OUTM CROSSP GND GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=2.4e+06u
X16_2 OUTM CROSSP GND GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=2.4e+06u
X17_0 OUTP CROSSN GND GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=2.4e+06u
X17_1 OUTP CROSSN GND GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=2.4e+06u
X17_2 OUTP CROSSN GND GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=2.4e+06u
X4_0 CROSSN CROSSP INTERN GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=2.4e+06u
X4_1 CROSSN CROSSP INTERN GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=2.4e+06u
X4_2 CROSSN CROSSP INTERN GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=2.4e+06u
X4_3 CROSSN CROSSP INTERN GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=2.4e+06u
X3_0 CROSSP CROSSN INTERP GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=2.4e+06u
X3_1 CROSSP CROSSN INTERP GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=2.4e+06u
X3_2 CROSSP CROSSN INTERP GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=2.4e+06u
X3_3 CROSSP CROSSN INTERP GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=2.4e+06u
X7_0 net050 CLK GND GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=2.16e+06u
X7_1 net050 CLK GND GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=2.16e+06u
X7_2 net050 CLK GND GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=2.16e+06u
X7_3 net050 CLK GND GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=2.16e+06u
X7_4 net050 CLK GND GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=2.16e+06u
X7_5 net050 CLK GND GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=2.16e+06u
X7_6 net050 CLK GND GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=2.16e+06u
X7_7 net050 CLK GND GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=2.16e+06u
X7_8 net050 CLK GND GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=2.16e+06u
X7_9 net050 CLK GND GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=2.16e+06u
X7_10 net050 CLK GND GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=2.16e+06u
X7_11 net050 CLK GND GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=2.16e+06u
X7_12 net050 CLK GND GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=2.16e+06u
X7_13 net050 CLK GND GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=2.16e+06u
X7_14 net050 CLK GND GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=2.16e+06u
X7_15 net050 CLK GND GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=2.16e+06u
X7_16 net050 CLK GND GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=2.16e+06u
X7_17 net050 CLK GND GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=2.16e+06u
X7_18 net050 CLK GND GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=2.16e+06u
X7_19 net050 CLK GND GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=2.16e+06u
X5_0 INTERN VI+ net050 GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=4.8e+06u
X5_1 INTERN VI+ net050 GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=4.8e+06u
X5_2 INTERN VI+ net050 GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=4.8e+06u
X5_3 INTERN VI+ net050 GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=4.8e+06u
X5_4 INTERN VI+ net050 GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=4.8e+06u
X5_5 INTERN VI+ net050 GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=4.8e+06u
X5_6 INTERN VI+ net050 GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=4.8e+06u
X5_7 INTERN VI+ net050 GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=4.8e+06u
X5_8 INTERN VI+ net050 GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=4.8e+06u
X5_9 INTERN VI+ net050 GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=4.8e+06u
X6_0 INTERP VI- net050 GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=4.8e+06u
X6_1 INTERP VI- net050 GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=4.8e+06u
X6_2 INTERP VI- net050 GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=4.8e+06u
X6_3 INTERP VI- net050 GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=4.8e+06u
X6_4 INTERP VI- net050 GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=4.8e+06u
X6_5 INTERP VI- net050 GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=4.8e+06u
X6_6 INTERP VI- net050 GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=4.8e+06u
X6_7 INTERP VI- net050 GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=4.8e+06u
X6_8 INTERP VI- net050 GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=4.8e+06u
X6_9 INTERP VI- net050 GND sky130_fd_pr__nfet_01v8_lvt l=2e+05u w=4.8e+06u
X8_0 OUTM CROSSP VDD VDD sky130_fd_pr__pfet_01v8 l=2e+05u w=4.8e+06u
X8_1 OUTM CROSSP VDD VDD sky130_fd_pr__pfet_01v8 l=2e+05u w=4.8e+06u
X8_2 OUTM CROSSP VDD VDD sky130_fd_pr__pfet_01v8 l=2e+05u w=4.8e+06u
X18_0 INTERN CLK VDD VDD sky130_fd_pr__pfet_01v8 l=2e+05u w=4.8e+06u
X18_1 INTERN CLK VDD VDD sky130_fd_pr__pfet_01v8 l=2e+05u w=4.8e+06u
X15_0 OUTP CROSSN VDD VDD sky130_fd_pr__pfet_01v8 l=2e+05u w=4.8e+06u
X15_1 OUTP CROSSN VDD VDD sky130_fd_pr__pfet_01v8 l=2e+05u w=4.8e+06u
X15_2 OUTP CROSSN VDD VDD sky130_fd_pr__pfet_01v8 l=2e+05u w=4.8e+06u
X19_0 INTERP CLK VDD VDD sky130_fd_pr__pfet_01v8 l=2e+05u w=4.8e+06u
X19_1 INTERP CLK VDD VDD sky130_fd_pr__pfet_01v8 l=2e+05u w=4.8e+06u
X10_0 CROSSN CLK VDD VDD sky130_fd_pr__pfet_01v8 l=2e+05u w=4.8e+06u
X10_1 CROSSN CLK VDD VDD sky130_fd_pr__pfet_01v8 l=2e+05u w=4.8e+06u
X12_0 CROSSP CLK VDD VDD sky130_fd_pr__pfet_01v8 l=2e+05u w=4.8e+06u
X12_1 CROSSP CLK VDD VDD sky130_fd_pr__pfet_01v8 l=2e+05u w=4.8e+06u
X14_0 CROSSN CROSSP VDD VDD sky130_fd_pr__pfet_01v8 l=2e+05u w=4.8e+06u
X14_1 CROSSN CROSSP VDD VDD sky130_fd_pr__pfet_01v8 l=2e+05u w=4.8e+06u
X14_2 CROSSN CROSSP VDD VDD sky130_fd_pr__pfet_01v8 l=2e+05u w=4.8e+06u
X14_3 CROSSN CROSSP VDD VDD sky130_fd_pr__pfet_01v8 l=2e+05u w=4.8e+06u
X13_0 CROSSP CROSSN VDD VDD sky130_fd_pr__pfet_01v8 l=2e+05u w=4.8e+06u
X13_1 CROSSP CROSSN VDD VDD sky130_fd_pr__pfet_01v8 l=2e+05u w=4.8e+06u
X13_2 CROSSP CROSSN VDD VDD sky130_fd_pr__pfet_01v8 l=2e+05u w=4.8e+06u
X13_3 CROSSP CROSSN VDD VDD sky130_fd_pr__pfet_01v8 l=2e+05u w=4.8e+06u

.ends
