VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  CAPACITANCE PICOFARADS 1 ;
  DATABASE MICRONS 2000 ;
END UNITS

MANUFACTURINGGRID 0.0005 ;

LAYER PO
  TYPE MASTERSLICE ;
END PO

LAYER CO
  TYPE CUT ;
END CO

LAYER M1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.52 0.52 ;
  WIDTH 0.14 ;
  AREA 0.083 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 
    WIDTH 0    0.14 
    WIDTH 3    0.28 ; 
END M1

LAYER VIA1
  TYPE CUT ;
  SPACING 0.17 ;
  WIDTH 0.15 ;
END VIA1

LAYER M2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.52 0.52 ;
  WIDTH 0.14 ;
  AREA 0.0676 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 
    WIDTH 0    0.14 
    WIDTH 3    0.28 ;
END M2

LAYER VIA2
  TYPE CUT ;
  SPACING 0.2 ;
  WIDTH 0.2 ;
END VIA2

LAYER M3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.36 0.36 ;
  WIDTH 0.3 ;
  AREA 0.24 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0
    WIDTH 0     0.3 
    WIDTH 3     0.4 ;
END M3

LAYER VIA3
  TYPE CUT ;
  SPACING 0.2 ;
  WIDTH 0.2 ;
END VIA3

LAYER M4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
  AREA 0.24 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0
    WIDTH 0     0.3 
    WIDTH 3     0.4 ;
END M4

LAYER VIA4
  TYPE CUT ;
  SPACING 0.8 ;
  WIDTH 0.8 ;
END VIA4

LAYER M5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
  AREA 0.4 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0
    WIDTH 0     1.6 ; 
END M5

VIARULE VIAG12 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.085 0.085 ;
    WIDTH 0.33 TO 4.50 ;
  LAYER M2 ;
    ENCLOSURE 0.085 0.085 ;
    WIDTH 0.33 TO 4.50 ;
  LAYER VIA1 ;
    RECT -0.075 -0.075 0.075 0.075 ;
    SPACING 0.32 BY 0.32 ;
END VIAG12

VIARULE VIAG23 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.085 0.085 ;
    WIDTH 0.33 TO 4.50 ;
  LAYER M3 ;
    ENCLOSURE 0.065 0.065 ;
    WIDTH 0.33 TO 4.50 ;
  LAYER VIA2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
    SPACING 0.4 BY 0.4 ;
END VIAG23

VIARULE VIAG34 GENERATE
  LAYER M3 ;
    ENCLOSURE 0.09 0.06 ;
    WIDTH 0.33 TO 4.50 ;
  LAYER M4 ;
    ENCLOSURE 0.065 0.065 ;
    WIDTH 0.33 TO 4.50 ;
  LAYER VIA2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
    SPACING 0.4 BY 0.4 ;
END VIAG34

VIARULE VIAG45 GENERATE
  LAYER M4 ;
    ENCLOSURE 0.19 0.19 ;
    WIDTH 0.33 TO 4.50 ;
  LAYER M5 ;
    ENCLOSURE 0.31 0.31 ;
    WIDTH 0.33 TO 4.50 ;
  LAYER VIA4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
    SPACING 1.6 BY 1.6 ;
END VIAG45

SITE CoreSite
  CLASS CORE ;
  SIZE 0.2 BY 1.71 ;
END CoreSite


END LIBRARY
