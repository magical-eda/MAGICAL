VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  CAPACITANCE PICOFARADS 1 ;
  DATABASE MICRONS 2000 ;
END UNITS

MANUFACTURINGGRID 0.0005 ;

LAYER PO
  TYPE MASTERSLICE ;
END PO

LAYER CO
  TYPE CUT ;
END CO

LAYER M1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.13 0.13 ;
  WIDTH 0.07 ;
  AREA 0.02 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 
    WIDTH 0    0.07 
    WIDTH 0.1  0.07 ; 
  SPACING 0.07 ENDOFLINE 0.07 WITHIN 0.025 ;
  MINSTEP 0.06 MAXEDGES 1 ;
END M1

LAYER VIA1
  TYPE CUT ;
  SPACING 0.07 ;
  WIDTH 0.07 ;
END VIA1

LAYER M2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.13 0.13 ;
  WIDTH 0.07 ;
  AREA 0.02 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 
    WIDTH 0    0.07 
    WIDTH 0.1  0.07 ;
  SPACING 0.07 ENDOFLINE 0.07 WITHIN 0.025 ;
  MINSTEP 0.06 MAXEDGES 1 ;
END M2

LAYER VIA2
  TYPE CUT ;
  SPACING 0.07 ;
  WIDTH 0.07 ;
END VIA2

LAYER M3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.13 0.13 ;
  WIDTH 0.07 ;
  AREA 0.02 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0
    WIDTH 0     0.07 
    WIDTH 0.1   0.07 ;
  SPACING 0.07 ENDOFLINE 0.07 WITHIN 0.035 ;
  MINSTEP 0.06 MAXEDGES 1 ;
END M3

LAYER VIA3
  TYPE CUT ;
  SPACING 0.07 ;
  WIDTH 0.07 ;
END VIA3

LAYER M4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.13 ;
  WIDTH 0.07 ;
  AREA 0.02 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0
    WIDTH 0     0.07 
    WIDTH 0.1   0.07 ;
  SPACING 0.07 ENDOFLINE 0.07 WITHIN 0.035 ;
  MINSTEP 0.06 MAXEDGES 1 ;
END M4

LAYER VIA4
  TYPE CUT ;
  SPACING 0.07 ;
  WIDTH 0.07 ;
END VIA4

LAYER M5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.13 ;
  WIDTH 0.07 ;
  AREA 0.02 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0
    WIDTH 0     0.07 
    WIDTH 0.1   0.07 ;
  SPACING 0.07 ENDOFLINE 0.07 WITHIN 0.035 ;
  MINSTEP 0.06 MAXEDGES 1 ;
END M5

LAYER VIA5
  TYPE CUT ;
  SPACING 0.07 ;
  WIDTH 0.07 ;
END VIA5

LAYER M6
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.13 ;
  WIDTH 0.07 ;
  AREA 0.02 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0
    WIDTH 0     0.07 
    WIDTH 0.1   0.07 ;
  SPACING 0.07 ENDOFLINE 0.07 WITHIN 0.035 ;
  MINSTEP 0.06 MAXEDGES 1 ;
END M6

LAYER VIA6
  TYPE CUT ;
  SPACING 0.07 ;
  WIDTH 0.07 ;
END VIA6

LAYER M7
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.13 ;
  WIDTH 0.07 ;
  AREA 0.02 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0
    WIDTH 0     0.07 
    WIDTH 0.1   0.07 ;
  SPACING 0.07 ENDOFLINE 0.07 WITHIN 0.035 ;
  MINSTEP 0.06 MAXEDGES 1 ;
END M7

VIA VIA12_1C DEFAULT 
    LAYER M1 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
    LAYER VIA1 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER M2 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA12_1C

VIA VIA12_1C_H DEFAULT 
    LAYER M1 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
    LAYER VIA1 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER M2 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA12_1C_H

VIA VIA12_1C_V DEFAULT 
    LAYER M1 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
    LAYER VIA1 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER M2 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA12_1C_V

VIA VIA23_1C DEFAULT 
    LAYER M2 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
    LAYER VIA2 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER M3 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA23_1C

VIA VIA23_1C_H DEFAULT 
    LAYER M2 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
    LAYER VIA2 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER M3 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA23_1C_H

VIA VIA23_1C_V DEFAULT 
    LAYER M2 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
    LAYER VIA2 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER M3 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA23_1C_V

VIA VIA23_1ST_N DEFAULT 
    LAYER M2 ;
        RECT -0.035000 -0.065000 0.035000 0.325000 ;
    LAYER VIA2 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER M3 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA23_1ST_N

VIA VIA23_1ST_S DEFAULT 
    LAYER M2 ;
        RECT -0.035000 -0.325000 0.035000 0.065000 ;
    LAYER VIA2 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER M3 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA23_1ST_S

VIA VIA34_1C DEFAULT 
    LAYER M3 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
    LAYER VIA3 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER M4 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA34_1C

VIA VIA34_1C_H DEFAULT 
    LAYER M3 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
    LAYER VIA3 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER M4 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA34_1C_H

VIA VIA34_1C_V DEFAULT 
    LAYER M3 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
    LAYER VIA3 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER M4 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA34_1C_V

VIA VIA34_1ST_E DEFAULT 
    LAYER M3 ;
        RECT -0.065000 -0.035000 0.325000 0.035000 ;
    LAYER VIA3 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER M4 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA34_1ST_E

VIA VIA34_1ST_W DEFAULT 
    LAYER M3 ;
        RECT -0.325000 -0.035000 0.065000 0.035000 ;
    LAYER VIA3 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER M4 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA34_1ST_W

VIA VIA45_1C DEFAULT 
    LAYER M4 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
    LAYER VIA4 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER M5 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA45_1C

VIA VIA45_1C_H DEFAULT 
    LAYER M4 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
    LAYER VIA4 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER M5 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA45_1C_H

VIA VIA45_1C_V DEFAULT 
    LAYER M4 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
    LAYER VIA4 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER M5 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA45_1C_V

VIA VIA45_1ST_N DEFAULT 
    LAYER M4 ;
        RECT -0.035000 -0.065000 0.035000 0.325000 ;
    LAYER VIA4 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER M5 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA45_1ST_N

VIA VIA45_1ST_S DEFAULT 
    LAYER M4 ;
        RECT -0.035000 -0.325000 0.035000 0.065000 ;
    LAYER VIA4 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER M5 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA45_1ST_S

VIA VIA5_0_VH DEFAULT 
    LAYER M5 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
    LAYER VIA5 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER M6 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA5_0_VH

VIA VIA6_0_HV DEFAULT 
    LAYER M6 ;
        RECT -0.260000 -0.200000 0.260000 0.200000 ;
    LAYER VIA6 ;
        RECT -0.180000 -0.180000 0.180000 0.180000 ;
    LAYER M7 ;
        RECT -0.200000 -0.260000 0.200000 0.260000 ;
END VIA6_0_HV


VIARULE VIAG12 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.03 0 ;
    WIDTH 0.10 TO 4.50 ;
  LAYER M2 ;
    ENCLOSURE 0.03 0 ;
    WIDTH 0.01 TO 4.50 ;
  LAYER VIA1 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.16 BY 0.16 ;
END VIAG12

VIARULE VIAG23 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.03 0 ;
    WIDTH 0.10 TO 4.50 ;
  LAYER M3 ;
    ENCLOSURE 0.03 0 ;
    WIDTH 0.01 TO 4.50 ;
  LAYER VIA2 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.16 BY 0.16 ;
END VIAG23

VIARULE VIAG34 GENERATE
  LAYER M3 ;
    ENCLOSURE 0.03 0 ;
    WIDTH 0.10 TO 4.50 ;
  LAYER M4 ;
    ENCLOSURE 0.03 0 ;
    WIDTH 0.01 TO 4.50 ;
  LAYER VIA2 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.16 BY 0.16 ;
END VIAG34

VIARULE VIAG45 GENERATE
  LAYER M4 ;
    ENCLOSURE 0.03 0 ;
    WIDTH 0.10 TO 4.50 ;
  LAYER M5 ;
    ENCLOSURE 0.03 0 ;
    WIDTH 0.01 TO 4.50 ;
  LAYER VIA4 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.16 BY 0.16 ;
END VIAG45

VIARULE VIAG56 GENERATE
  LAYER M5 ;
    ENCLOSURE 0.03 0 ;
    WIDTH 0.10 TO 4.50 ;
  LAYER M6 ;
    ENCLOSURE 0.03 0 ;
    WIDTH 0.01 TO 4.50 ;
  LAYER VIA5 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.16 BY 0.16 ;
END VIAG56

VIARULE VIAG67 GENERATE
  LAYER M6 ;
    ENCLOSURE 0.03 0 ;
    WIDTH 0.10 TO 4.50 ;
  LAYER M7 ;
    ENCLOSURE 0.03 0 ;
    WIDTH 0.01 TO 4.50 ;
  LAYER VIA6 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.16 BY 0.16 ;
END VIAG67


SITE CoreSite
  CLASS CORE ;
  SIZE 0.2 BY 1.71 ;
END CoreSite


END LIBRARY
